library verilog;
use verilog.vl_types.all;
entity TB_contadorMod16 is
end TB_contadorMod16;
