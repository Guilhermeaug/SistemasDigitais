library verilog;
use verilog.vl_types.all;
entity TB_contadorMod13 is
end TB_contadorMod13;
